library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package ram_data_width_pkg is

    constant ram_port_width : integer := 16;

end package ram_data_width_pkg;
------------------------------------------------------------------------
